//`include "axi_interface.sv"

package axi_pkg;
`include "uvm_macros.svh"
import uvm_pkg::*;
import cmd_pkg::*;

`include "axi_config.sv"
`include "valid_data.sv"
`include "hmc_pkt_item_request.sv"
`include "axi_sequencer.sv"
`include "axi_driver.sv"
`include "axi_monitor.sv"
`include "axi_agent.sv" 


endpackage : axi_pkg
