package rf_reg_block_pkg;
  
  //uvm pakage and macros
  import uvm_pkg::*;
  `include "uvm_macros.svh"


`include "reg_error_abort_not_cleared.sv"
`include "reg_counter_reset.sv"
`include "reg_errors_on_rx.sv"
`include "reg_poisoned_packets.sv"
`include "reg_rcvd_rsp.sv"
`include "reg_run_length_bit_flip.sv"
`include "reg_sent_np.sv"
`include "reg_sent_p.sv"
`include "reg_sent_r.sv"
`include "reg_status_general.sv"
`include "reg_status_init.sv"
`include "reg_tx_link_retries.sv"
`include "reg_control.sv"

`include "rf_reg_block.sv"
  
endpackage : rf_reg_block_pkg